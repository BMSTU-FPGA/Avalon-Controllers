
module TEST_OY_CPU (
	clk_clk,
	mealymoure_mm_controller_0_ledg_export,
	mealymoure_mm_controller_0_ledr_export);	

	input		clk_clk;
	output	[8:0]	mealymoure_mm_controller_0_ledg_export;
	output	[17:0]	mealymoure_mm_controller_0_ledr_export;
endmodule
