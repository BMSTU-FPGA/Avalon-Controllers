-- TEST_OY_CPU.vhd

-- Generated using ACDS version 23.1 993

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity TEST_OY_CPU is
	port (
		clk_clk : in std_logic := '0'  -- clk.clk
	);
end entity TEST_OY_CPU;

architecture rtl of TEST_OY_CPU is
	component Number_generator_controller is
		port (
			avs_s0_chipselect : in  std_logic                     := 'X';             -- chipselect
			avs_s0_byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avs_s0_read       : in  std_logic                     := 'X';             -- read
			avs_s0_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			avs_s0_write      : in  std_logic                     := 'X';             -- write
			avs_s0_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			csi_clk           : in  std_logic                     := 'X';             -- clk
			rsi_reset         : in  std_logic                     := 'X'              -- reset
		);
	end component Number_generator_controller;

	component CI_NG is
		port (
			clk    : in  std_logic                     := 'X'; -- clk
			result : out std_logic_vector(31 downto 0);        -- result
			resetn : in  std_logic                     := 'X'  -- reset_n
		);
	end component CI_NG;

	component OY_Instruction_Controller is
		generic (
			n : integer := 16
		);
		port (
			ncs_clk    : in  std_logic                     := 'X';             -- clk
			ncs_reset  : in  std_logic                     := 'X';             -- reset
			ncs_start  : in  std_logic                     := 'X';             -- start
			ncs_dataa  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ncs_datab  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ncs_done   : out std_logic;                                        -- done
			ncs_result : out std_logic_vector(31 downto 0)                     -- result
		);
	end component OY_Instruction_Controller;

	component OY_MM_Controller is
		generic (
			n : integer := 16
		);
		port (
			avs_chipselect  : in  std_logic                     := 'X';             -- chipselect
			avs_address     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			avs_read        : in  std_logic                     := 'X';             -- read
			avs_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			avs_write       : in  std_logic                     := 'X';             -- write
			avs_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avs_waitrequest : out std_logic;                                        -- waitrequest
			csi_clk         : in  std_logic                     := 'X';             -- clk
			rsi_reset       : in  std_logic                     := 'X';             -- reset
			ins_irq         : out std_logic                                         -- irq
		);
	end component OY_MM_Controller;

	component TEST_OY_Controller is
		generic (
			n : integer := 16
		);
		port (
			avs_chipselect  : in  std_logic                     := 'X';             -- chipselect
			avs_address     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			avs_read        : in  std_logic                     := 'X';             -- read
			avs_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			avs_write       : in  std_logic                     := 'X';             -- write
			avs_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avs_waitrequest : out std_logic;                                        -- waitrequest
			csi_clk         : in  std_logic                     := 'X';             -- clk
			rsi_reset       : in  std_logic                     := 'X';             -- reset
			ins_irq         : out std_logic                                         -- irq
		);
	end component TEST_OY_Controller;

	component TEST_OY_CPU_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(13 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(13 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			E_ci_multi_done                     : in  std_logic                     := 'X';             -- done
			E_ci_multi_clk_en                   : out std_logic;                                        -- clk_en
			E_ci_multi_start                    : out std_logic;                                        -- start
			E_ci_result                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			D_ci_a                              : out std_logic_vector(4 downto 0);                     -- a
			D_ci_b                              : out std_logic_vector(4 downto 0);                     -- b
			D_ci_c                              : out std_logic_vector(4 downto 0);                     -- c
			D_ci_n                              : out std_logic_vector(7 downto 0);                     -- n
			D_ci_readra                         : out std_logic;                                        -- readra
			D_ci_readrb                         : out std_logic;                                        -- readrb
			D_ci_writerc                        : out std_logic;                                        -- writerc
			E_ci_dataa                          : out std_logic_vector(31 downto 0);                    -- dataa
			E_ci_datab                          : out std_logic_vector(31 downto 0);                    -- datab
			E_ci_multi_clock                    : out std_logic;                                        -- clk
			E_ci_multi_reset                    : out std_logic;                                        -- reset
			E_ci_multi_reset_req                : out std_logic;                                        -- reset_req
			W_ci_estatus                        : out std_logic;                                        -- estatus
			W_ci_ipending                       : out std_logic_vector(31 downto 0)                     -- ipending
		);
	end component TEST_OY_CPU_nios2_gen2_0;

	component TEST_OY_CPU_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component TEST_OY_CPU_onchip_memory2_0;

	component altera_customins_master_translator is
		generic (
			SHARED_COMB_AND_MULTI : integer := 0
		);
		port (
			ci_slave_dataa            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result           : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n                : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra           : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb           : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc          : in  std_logic                     := 'X';             -- writerc
			ci_slave_a                : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b                : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c                : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus          : in  std_logic                     := 'X';             -- estatus
			ci_slave_multi_clk        : in  std_logic                     := 'X';             -- clk
			ci_slave_multi_reset      : in  std_logic                     := 'X';             -- reset
			ci_slave_multi_clken      : in  std_logic                     := 'X';             -- clk_en
			ci_slave_multi_reset_req  : in  std_logic                     := 'X';             -- reset_req
			ci_slave_multi_start      : in  std_logic                     := 'X';             -- start
			ci_slave_multi_done       : out std_logic;                                        -- done
			comb_ci_master_dataa      : out std_logic_vector(31 downto 0);                    -- dataa
			comb_ci_master_datab      : out std_logic_vector(31 downto 0);                    -- datab
			comb_ci_master_result     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			comb_ci_master_n          : out std_logic_vector(7 downto 0);                     -- n
			comb_ci_master_readra     : out std_logic;                                        -- readra
			comb_ci_master_readrb     : out std_logic;                                        -- readrb
			comb_ci_master_writerc    : out std_logic;                                        -- writerc
			comb_ci_master_a          : out std_logic_vector(4 downto 0);                     -- a
			comb_ci_master_b          : out std_logic_vector(4 downto 0);                     -- b
			comb_ci_master_c          : out std_logic_vector(4 downto 0);                     -- c
			comb_ci_master_ipending   : out std_logic_vector(31 downto 0);                    -- ipending
			comb_ci_master_estatus    : out std_logic;                                        -- estatus
			multi_ci_master_clk       : out std_logic;                                        -- clk
			multi_ci_master_reset     : out std_logic;                                        -- reset
			multi_ci_master_clken     : out std_logic;                                        -- clk_en
			multi_ci_master_reset_req : out std_logic;                                        -- reset_req
			multi_ci_master_start     : out std_logic;                                        -- start
			multi_ci_master_done      : in  std_logic                     := 'X';             -- done
			multi_ci_master_dataa     : out std_logic_vector(31 downto 0);                    -- dataa
			multi_ci_master_datab     : out std_logic_vector(31 downto 0);                    -- datab
			multi_ci_master_result    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			multi_ci_master_n         : out std_logic_vector(7 downto 0);                     -- n
			multi_ci_master_readra    : out std_logic;                                        -- readra
			multi_ci_master_readrb    : out std_logic;                                        -- readrb
			multi_ci_master_writerc   : out std_logic;                                        -- writerc
			multi_ci_master_a         : out std_logic_vector(4 downto 0);                     -- a
			multi_ci_master_b         : out std_logic_vector(4 downto 0);                     -- b
			multi_ci_master_c         : out std_logic_vector(4 downto 0);                     -- c
			ci_slave_multi_dataa      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_dataa
			ci_slave_multi_datab      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_datab
			ci_slave_multi_result     : out std_logic_vector(31 downto 0);                    -- multi_result
			ci_slave_multi_n          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- multi_n
			ci_slave_multi_readra     : in  std_logic                     := 'X';             -- multi_readra
			ci_slave_multi_readrb     : in  std_logic                     := 'X';             -- multi_readrb
			ci_slave_multi_writerc    : in  std_logic                     := 'X';             -- multi_writerc
			ci_slave_multi_a          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_a
			ci_slave_multi_b          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_b
			ci_slave_multi_c          : in  std_logic_vector(4 downto 0)  := (others => 'X')  -- multi_c
		);
	end component altera_customins_master_translator;

	component TEST_OY_CPU_nios2_gen2_0_custom_instruction_master_comb_xconnect is
		port (
			ci_slave_dataa      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result     : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra     : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb     : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc    : in  std_logic                     := 'X';             -- writerc
			ci_slave_a          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus    : in  std_logic                     := 'X';             -- estatus
			ci_master0_dataa    : out std_logic_vector(31 downto 0);                    -- dataa
			ci_master0_datab    : out std_logic_vector(31 downto 0);                    -- datab
			ci_master0_result   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			ci_master0_n        : out std_logic_vector(7 downto 0);                     -- n
			ci_master0_readra   : out std_logic;                                        -- readra
			ci_master0_readrb   : out std_logic;                                        -- readrb
			ci_master0_writerc  : out std_logic;                                        -- writerc
			ci_master0_a        : out std_logic_vector(4 downto 0);                     -- a
			ci_master0_b        : out std_logic_vector(4 downto 0);                     -- b
			ci_master0_c        : out std_logic_vector(4 downto 0);                     -- c
			ci_master0_ipending : out std_logic_vector(31 downto 0);                    -- ipending
			ci_master0_estatus  : out std_logic                                         -- estatus
		);
	end component TEST_OY_CPU_nios2_gen2_0_custom_instruction_master_comb_xconnect;

	component TEST_OY_CPU_nios2_gen2_0_custom_instruction_master_multi_xconnect is
		port (
			ci_slave_dataa       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result      : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra      : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb      : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc     : in  std_logic                     := 'X';             -- writerc
			ci_slave_a           : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b           : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c           : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus     : in  std_logic                     := 'X';             -- estatus
			ci_slave_clk         : in  std_logic                     := 'X';             -- clk
			ci_slave_reset       : in  std_logic                     := 'X';             -- reset
			ci_slave_clken       : in  std_logic                     := 'X';             -- clk_en
			ci_slave_reset_req   : in  std_logic                     := 'X';             -- reset_req
			ci_slave_start       : in  std_logic                     := 'X';             -- start
			ci_slave_done        : out std_logic;                                        -- done
			ci_master0_dataa     : out std_logic_vector(31 downto 0);                    -- dataa
			ci_master0_datab     : out std_logic_vector(31 downto 0);                    -- datab
			ci_master0_result    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			ci_master0_n         : out std_logic_vector(7 downto 0);                     -- n
			ci_master0_readra    : out std_logic;                                        -- readra
			ci_master0_readrb    : out std_logic;                                        -- readrb
			ci_master0_writerc   : out std_logic;                                        -- writerc
			ci_master0_a         : out std_logic_vector(4 downto 0);                     -- a
			ci_master0_b         : out std_logic_vector(4 downto 0);                     -- b
			ci_master0_c         : out std_logic_vector(4 downto 0);                     -- c
			ci_master0_ipending  : out std_logic_vector(31 downto 0);                    -- ipending
			ci_master0_estatus   : out std_logic;                                        -- estatus
			ci_master0_clk       : out std_logic;                                        -- clk
			ci_master0_reset     : out std_logic;                                        -- reset
			ci_master0_clken     : out std_logic;                                        -- clk_en
			ci_master0_reset_req : out std_logic;                                        -- reset_req
			ci_master0_start     : out std_logic;                                        -- start
			ci_master0_done      : in  std_logic                     := 'X'              -- done
		);
	end component TEST_OY_CPU_nios2_gen2_0_custom_instruction_master_multi_xconnect;

	component TEST_OY_CPU_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                        : in  std_logic                     := 'X';             -- clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset       : in  std_logic                     := 'X';             -- reset
			OY_MM_Controller_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address                     : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest                 : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable                  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                        : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata                    : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_write                       : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess                 : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest          : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read                 : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			NG_Controller_0_s0_write                             : out std_logic;                                        -- write
			NG_Controller_0_s0_read                              : out std_logic;                                        -- read
			NG_Controller_0_s0_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			NG_Controller_0_s0_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			NG_Controller_0_s0_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			NG_Controller_0_s0_chipselect                        : out std_logic;                                        -- chipselect
			nios2_gen2_0_debug_mem_slave_address                 : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write                   : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read                    : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable              : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest             : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess             : out std_logic;                                        -- debugaccess
			onchip_memory2_0_s1_address                          : out std_logic_vector(9 downto 0);                     -- address
			onchip_memory2_0_s1_write                            : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                       : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                       : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                            : out std_logic;                                        -- clken
			OY_MM_Controller_0_avalon_slave_0_address            : out std_logic_vector(1 downto 0);                     -- address
			OY_MM_Controller_0_avalon_slave_0_write              : out std_logic;                                        -- write
			OY_MM_Controller_0_avalon_slave_0_read               : out std_logic;                                        -- read
			OY_MM_Controller_0_avalon_slave_0_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			OY_MM_Controller_0_avalon_slave_0_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			OY_MM_Controller_0_avalon_slave_0_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			OY_MM_Controller_0_avalon_slave_0_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			OY_MM_Controller_0_avalon_slave_0_chipselect         : out std_logic;                                        -- chipselect
			TEST_OY_Controller_0_avalon_slave_0_address          : out std_logic_vector(1 downto 0);                     -- address
			TEST_OY_Controller_0_avalon_slave_0_write            : out std_logic;                                        -- write
			TEST_OY_Controller_0_avalon_slave_0_read             : out std_logic;                                        -- read
			TEST_OY_Controller_0_avalon_slave_0_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TEST_OY_Controller_0_avalon_slave_0_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			TEST_OY_Controller_0_avalon_slave_0_byteenable       : out std_logic_vector(3 downto 0);                     -- byteenable
			TEST_OY_Controller_0_avalon_slave_0_waitrequest      : in  std_logic                     := 'X';             -- waitrequest
			TEST_OY_Controller_0_avalon_slave_0_chipselect       : out std_logic                                         -- chipselect
		);
	end component TEST_OY_CPU_mm_interconnect_0;

	component TEST_OY_CPU_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component TEST_OY_CPU_irq_mapper;

	component test_oy_cpu_nios2_gen2_0_custom_instruction_master_comb_slave_translator0 is
		generic (
			N_WIDTH          : integer := 8;
			USE_DONE         : integer := 1;
			NUM_FIXED_CYCLES : integer := 2
		);
		port (
			ci_slave_dataa      : in  std_logic_vector(31 downto 0) := (others => 'X'); --  ci_slave.dataa
			ci_slave_datab      : in  std_logic_vector(31 downto 0) := (others => 'X'); --          .datab
			ci_slave_result     : out std_logic_vector(31 downto 0);                    --          .result
			ci_slave_n          : in  std_logic_vector(7 downto 0)  := (others => 'X'); --          .n
			ci_slave_readra     : in  std_logic                     := 'X';             --          .readra
			ci_slave_readrb     : in  std_logic                     := 'X';             --          .readrb
			ci_slave_writerc    : in  std_logic                     := 'X';             --          .writerc
			ci_slave_a          : in  std_logic_vector(4 downto 0)  := (others => 'X'); --          .a
			ci_slave_b          : in  std_logic_vector(4 downto 0)  := (others => 'X'); --          .b
			ci_slave_c          : in  std_logic_vector(4 downto 0)  := (others => 'X'); --          .c
			ci_slave_ipending   : in  std_logic_vector(31 downto 0) := (others => 'X'); --          .ipending
			ci_slave_estatus    : in  std_logic                     := 'X';             --          .estatus
			ci_master_result    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ci_master.result
			ci_master_a         : out std_logic_vector(4 downto 0);
			ci_master_b         : out std_logic_vector(4 downto 0);
			ci_master_c         : out std_logic_vector(4 downto 0);
			ci_master_clk       : out std_logic;
			ci_master_clken     : out std_logic;
			ci_master_dataa     : out std_logic_vector(31 downto 0);
			ci_master_datab     : out std_logic_vector(31 downto 0);
			ci_master_done      : in  std_logic                     := 'X';
			ci_master_estatus   : out std_logic;
			ci_master_ipending  : out std_logic_vector(31 downto 0);
			ci_master_n         : out std_logic_vector(7 downto 0);
			ci_master_readra    : out std_logic;
			ci_master_readrb    : out std_logic;
			ci_master_reset     : out std_logic;
			ci_master_reset_req : out std_logic;
			ci_master_start     : out std_logic;
			ci_master_writerc   : out std_logic;
			ci_slave_clk        : in  std_logic                     := 'X';
			ci_slave_clken      : in  std_logic                     := 'X';
			ci_slave_done       : out std_logic;
			ci_slave_reset      : in  std_logic                     := 'X';
			ci_slave_reset_req  : in  std_logic                     := 'X';
			ci_slave_start      : in  std_logic                     := 'X'
		);
	end component test_oy_cpu_nios2_gen2_0_custom_instruction_master_comb_slave_translator0;

	component test_oy_cpu_nios2_gen2_0_custom_instruction_master_multi_slave_translator0 is
		generic (
			N_WIDTH          : integer := 8;
			USE_DONE         : integer := 1;
			NUM_FIXED_CYCLES : integer := 2
		);
		port (
			ci_slave_dataa      : in  std_logic_vector(31 downto 0) := (others => 'X'); --  ci_slave.dataa
			ci_slave_datab      : in  std_logic_vector(31 downto 0) := (others => 'X'); --          .datab
			ci_slave_result     : out std_logic_vector(31 downto 0);                    --          .result
			ci_slave_n          : in  std_logic_vector(7 downto 0)  := (others => 'X'); --          .n
			ci_slave_readra     : in  std_logic                     := 'X';             --          .readra
			ci_slave_readrb     : in  std_logic                     := 'X';             --          .readrb
			ci_slave_writerc    : in  std_logic                     := 'X';             --          .writerc
			ci_slave_a          : in  std_logic_vector(4 downto 0)  := (others => 'X'); --          .a
			ci_slave_b          : in  std_logic_vector(4 downto 0)  := (others => 'X'); --          .b
			ci_slave_c          : in  std_logic_vector(4 downto 0)  := (others => 'X'); --          .c
			ci_slave_ipending   : in  std_logic_vector(31 downto 0) := (others => 'X'); --          .ipending
			ci_slave_estatus    : in  std_logic                     := 'X';             --          .estatus
			ci_slave_clk        : in  std_logic                     := 'X';             --          .clk
			ci_slave_clken      : in  std_logic                     := 'X';             --          .clk_en
			ci_slave_reset_req  : in  std_logic                     := 'X';             --          .reset_req
			ci_slave_reset      : in  std_logic                     := 'X';             --          .reset
			ci_slave_start      : in  std_logic                     := 'X';             --          .start
			ci_slave_done       : out std_logic;                                        --          .done
			ci_master_dataa     : out std_logic_vector(31 downto 0);                    -- ci_master.dataa
			ci_master_datab     : out std_logic_vector(31 downto 0);                    --          .datab
			ci_master_result    : in  std_logic_vector(31 downto 0) := (others => 'X'); --          .result
			ci_master_clk       : out std_logic;                                        --          .clk
			ci_master_clken     : out std_logic;                                        --          .clk_en
			ci_master_reset     : out std_logic;                                        --          .reset
			ci_master_start     : out std_logic;                                        --          .start
			ci_master_done      : in  std_logic                     := 'X';             --          .done
			ci_master_a         : out std_logic_vector(4 downto 0);
			ci_master_b         : out std_logic_vector(4 downto 0);
			ci_master_c         : out std_logic_vector(4 downto 0);
			ci_master_estatus   : out std_logic;
			ci_master_ipending  : out std_logic_vector(31 downto 0);
			ci_master_n         : out std_logic_vector(7 downto 0);
			ci_master_readra    : out std_logic;
			ci_master_readrb    : out std_logic;
			ci_master_reset_req : out std_logic;
			ci_master_writerc   : out std_logic
		);
	end component test_oy_cpu_nios2_gen2_0_custom_instruction_master_multi_slave_translator0;

	component test_oy_cpu_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component test_oy_cpu_rst_controller;

	component test_oy_cpu_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component test_oy_cpu_rst_controller_001;

	signal nios2_gen2_0_debug_reset_request_reset                                          : std_logic;                     -- nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in0, rst_controller:reset_in1, rst_controller_001:reset_in0]
	signal nios2_gen2_0_custom_instruction_master_readra                                   : std_logic;                     -- nios2_gen2_0:D_ci_readra -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_readra
	signal nios2_gen2_0_custom_instruction_master_a                                        : std_logic_vector(4 downto 0);  -- nios2_gen2_0:D_ci_a -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_a
	signal nios2_gen2_0_custom_instruction_master_b                                        : std_logic_vector(4 downto 0);  -- nios2_gen2_0:D_ci_b -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_b
	signal nios2_gen2_0_custom_instruction_master_c                                        : std_logic_vector(4 downto 0);  -- nios2_gen2_0:D_ci_c -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_c
	signal nios2_gen2_0_custom_instruction_master_readrb                                   : std_logic;                     -- nios2_gen2_0:D_ci_readrb -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_readrb
	signal nios2_gen2_0_custom_instruction_master_clk                                      : std_logic;                     -- nios2_gen2_0:E_ci_multi_clock -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_clk
	signal nios2_gen2_0_custom_instruction_master_ipending                                 : std_logic_vector(31 downto 0); -- nios2_gen2_0:W_ci_ipending -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_ipending
	signal nios2_gen2_0_custom_instruction_master_start                                    : std_logic;                     -- nios2_gen2_0:E_ci_multi_start -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_start
	signal nios2_gen2_0_custom_instruction_master_reset_req                                : std_logic;                     -- nios2_gen2_0:E_ci_multi_reset_req -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_reset_req
	signal nios2_gen2_0_custom_instruction_master_done                                     : std_logic;                     -- nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_done -> nios2_gen2_0:E_ci_multi_done
	signal nios2_gen2_0_custom_instruction_master_n                                        : std_logic_vector(7 downto 0);  -- nios2_gen2_0:D_ci_n -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_n
	signal nios2_gen2_0_custom_instruction_master_result                                   : std_logic_vector(31 downto 0); -- nios2_gen2_0_custom_instruction_master_translator:ci_slave_result -> nios2_gen2_0:E_ci_result
	signal nios2_gen2_0_custom_instruction_master_estatus                                  : std_logic;                     -- nios2_gen2_0:W_ci_estatus -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_estatus
	signal nios2_gen2_0_custom_instruction_master_clk_en                                   : std_logic;                     -- nios2_gen2_0:E_ci_multi_clk_en -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_clken
	signal nios2_gen2_0_custom_instruction_master_datab                                    : std_logic_vector(31 downto 0); -- nios2_gen2_0:E_ci_datab -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_datab
	signal nios2_gen2_0_custom_instruction_master_dataa                                    : std_logic_vector(31 downto 0); -- nios2_gen2_0:E_ci_dataa -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_dataa
	signal nios2_gen2_0_custom_instruction_master_reset                                    : std_logic;                     -- nios2_gen2_0:E_ci_multi_reset -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_reset
	signal nios2_gen2_0_custom_instruction_master_writerc                                  : std_logic;                     -- nios2_gen2_0:D_ci_writerc -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_writerc
	signal nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_result         : std_logic_vector(31 downto 0); -- nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_result -> nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_result
	signal nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_readra         : std_logic;                     -- nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_readra -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_readra
	signal nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_a              : std_logic_vector(4 downto 0);  -- nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_a -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_a
	signal nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_b              : std_logic_vector(4 downto 0);  -- nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_b -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_b
	signal nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_readrb         : std_logic;                     -- nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_readrb -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_readrb
	signal nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_c              : std_logic_vector(4 downto 0);  -- nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_c -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_c
	signal nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_estatus        : std_logic;                     -- nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_estatus -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_estatus
	signal nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_ipending       : std_logic_vector(31 downto 0); -- nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_ipending -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_ipending
	signal nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_datab          : std_logic_vector(31 downto 0); -- nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_datab -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_datab
	signal nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_dataa          : std_logic_vector(31 downto 0); -- nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_dataa -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_dataa
	signal nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_writerc        : std_logic;                     -- nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_writerc -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_writerc
	signal nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_n              : std_logic_vector(7 downto 0);  -- nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_n -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_n
	signal nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_result          : std_logic_vector(31 downto 0); -- nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_result -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_result
	signal nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_readra          : std_logic;                     -- nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_readra -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	signal nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_a               : std_logic_vector(4 downto 0);  -- nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_a -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_a
	signal nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_b               : std_logic_vector(4 downto 0);  -- nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_b -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_b
	signal nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_readrb          : std_logic;                     -- nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_readrb -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	signal nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_c               : std_logic_vector(4 downto 0);  -- nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_c -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_c
	signal nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_estatus         : std_logic;                     -- nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_estatus -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	signal nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_ipending        : std_logic_vector(31 downto 0); -- nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_ipending -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	signal nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_datab           : std_logic_vector(31 downto 0); -- nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_datab -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	signal nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_dataa           : std_logic_vector(31 downto 0); -- nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_dataa -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	signal nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_writerc         : std_logic;                     -- nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_writerc -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	signal nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_n               : std_logic_vector(7 downto 0);  -- nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_n -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_n
	signal nios2_gen2_0_custom_instruction_master_comb_slave_translator0_ci_master_result  : std_logic_vector(31 downto 0); -- NG_Instr_Controller_0:result -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_master_result
	signal nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_readra        : std_logic;                     -- nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_readra -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_readra
	signal nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_a             : std_logic_vector(4 downto 0);  -- nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_a -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_a
	signal nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_b             : std_logic_vector(4 downto 0);  -- nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_b -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_b
	signal nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_clk           : std_logic;                     -- nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_clk -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_clk
	signal nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_readrb        : std_logic;                     -- nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_readrb -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_readrb
	signal nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_c             : std_logic_vector(4 downto 0);  -- nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_c -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_c
	signal nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_start         : std_logic;                     -- nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_start -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_start
	signal nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_reset_req     : std_logic;                     -- nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_reset_req -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	signal nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_done          : std_logic;                     -- nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_done -> nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_done
	signal nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_n             : std_logic_vector(7 downto 0);  -- nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_n -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_n
	signal nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_result        : std_logic_vector(31 downto 0); -- nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_result -> nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_result
	signal nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_clk_en        : std_logic;                     -- nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_clken -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_clken
	signal nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_datab         : std_logic_vector(31 downto 0); -- nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_datab -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_datab
	signal nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_dataa         : std_logic_vector(31 downto 0); -- nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_dataa -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_dataa
	signal nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_reset         : std_logic;                     -- nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_reset -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_reset
	signal nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_writerc       : std_logic;                     -- nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_writerc -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_writerc
	signal nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_readra         : std_logic;                     -- nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_readra -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	signal nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_a              : std_logic_vector(4 downto 0);  -- nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_a -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_a
	signal nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_b              : std_logic_vector(4 downto 0);  -- nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_b -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_b
	signal nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_readrb         : std_logic;                     -- nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_readrb -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	signal nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_c              : std_logic_vector(4 downto 0);  -- nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_c -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_c
	signal nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_clk            : std_logic;                     -- nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_clk -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	signal nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_ipending       : std_logic_vector(31 downto 0); -- nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_ipending -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	signal nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_start          : std_logic;                     -- nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_start -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_start
	signal nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_reset_req      : std_logic;                     -- nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	signal nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_done           : std_logic;                     -- nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_done -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_done
	signal nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_n              : std_logic_vector(7 downto 0);  -- nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_n -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_n
	signal nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_result         : std_logic_vector(31 downto 0); -- nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_result -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_result
	signal nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_estatus        : std_logic;                     -- nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_estatus -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	signal nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_clk_en         : std_logic;                     -- nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_clken -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	signal nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_datab          : std_logic_vector(31 downto 0); -- nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_datab -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	signal nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_dataa          : std_logic_vector(31 downto 0); -- nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_dataa -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	signal nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_reset          : std_logic;                     -- nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_reset -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	signal nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_writerc        : std_logic;                     -- nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_writerc -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	signal nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_result : std_logic_vector(31 downto 0); -- OY_Instr_Controller_0:ncs_result -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_result
	signal nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_clk    : std_logic;                     -- nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_clk -> OY_Instr_Controller_0:ncs_clk
	signal nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_datab  : std_logic_vector(31 downto 0); -- nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_datab -> OY_Instr_Controller_0:ncs_datab
	signal nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_dataa  : std_logic_vector(31 downto 0); -- nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> OY_Instr_Controller_0:ncs_dataa
	signal nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_start  : std_logic;                     -- nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_start -> OY_Instr_Controller_0:ncs_start
	signal nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_reset  : std_logic;                     -- nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_reset -> OY_Instr_Controller_0:ncs_reset
	signal nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_done   : std_logic;                     -- OY_Instr_Controller_0:ncs_done -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_done
	signal nios2_gen2_0_data_master_readdata                                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                                            : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                                            : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                                : std_logic_vector(13 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                                             : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                                   : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                                                  : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                                              : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                                     : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                                         : std_logic_vector(13 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                                            : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_chipselect                  : std_logic;                     -- mm_interconnect_0:OY_MM_Controller_0_avalon_slave_0_chipselect -> OY_MM_Controller_0:avs_chipselect
	signal mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_readdata                    : std_logic_vector(31 downto 0); -- OY_MM_Controller_0:avs_readdata -> mm_interconnect_0:OY_MM_Controller_0_avalon_slave_0_readdata
	signal mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_waitrequest                 : std_logic;                     -- OY_MM_Controller_0:avs_waitrequest -> mm_interconnect_0:OY_MM_Controller_0_avalon_slave_0_waitrequest
	signal mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_address                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:OY_MM_Controller_0_avalon_slave_0_address -> OY_MM_Controller_0:avs_address
	signal mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_read                        : std_logic;                     -- mm_interconnect_0:OY_MM_Controller_0_avalon_slave_0_read -> OY_MM_Controller_0:avs_read
	signal mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_byteenable                  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:OY_MM_Controller_0_avalon_slave_0_byteenable -> OY_MM_Controller_0:avs_byteenable
	signal mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_write                       : std_logic;                     -- mm_interconnect_0:OY_MM_Controller_0_avalon_slave_0_write -> OY_MM_Controller_0:avs_write
	signal mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:OY_MM_Controller_0_avalon_slave_0_writedata -> OY_MM_Controller_0:avs_writedata
	signal mm_interconnect_0_test_oy_controller_0_avalon_slave_0_chipselect                : std_logic;                     -- mm_interconnect_0:TEST_OY_Controller_0_avalon_slave_0_chipselect -> TEST_OY_Controller_0:avs_chipselect
	signal mm_interconnect_0_test_oy_controller_0_avalon_slave_0_readdata                  : std_logic_vector(31 downto 0); -- TEST_OY_Controller_0:avs_readdata -> mm_interconnect_0:TEST_OY_Controller_0_avalon_slave_0_readdata
	signal mm_interconnect_0_test_oy_controller_0_avalon_slave_0_waitrequest               : std_logic;                     -- TEST_OY_Controller_0:avs_waitrequest -> mm_interconnect_0:TEST_OY_Controller_0_avalon_slave_0_waitrequest
	signal mm_interconnect_0_test_oy_controller_0_avalon_slave_0_address                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:TEST_OY_Controller_0_avalon_slave_0_address -> TEST_OY_Controller_0:avs_address
	signal mm_interconnect_0_test_oy_controller_0_avalon_slave_0_read                      : std_logic;                     -- mm_interconnect_0:TEST_OY_Controller_0_avalon_slave_0_read -> TEST_OY_Controller_0:avs_read
	signal mm_interconnect_0_test_oy_controller_0_avalon_slave_0_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:TEST_OY_Controller_0_avalon_slave_0_byteenable -> TEST_OY_Controller_0:avs_byteenable
	signal mm_interconnect_0_test_oy_controller_0_avalon_slave_0_write                     : std_logic;                     -- mm_interconnect_0:TEST_OY_Controller_0_avalon_slave_0_write -> TEST_OY_Controller_0:avs_write
	signal mm_interconnect_0_test_oy_controller_0_avalon_slave_0_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:TEST_OY_Controller_0_avalon_slave_0_writedata -> TEST_OY_Controller_0:avs_writedata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata                         : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest                      : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess                      : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address                          : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read                             : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable                       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write                            : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_ng_controller_0_s0_chipselect                                 : std_logic;                     -- mm_interconnect_0:NG_Controller_0_s0_chipselect -> NG_Controller_0:avs_s0_chipselect
	signal mm_interconnect_0_ng_controller_0_s0_readdata                                   : std_logic_vector(31 downto 0); -- NG_Controller_0:avs_s0_readdata -> mm_interconnect_0:NG_Controller_0_s0_readdata
	signal mm_interconnect_0_ng_controller_0_s0_read                                       : std_logic;                     -- mm_interconnect_0:NG_Controller_0_s0_read -> NG_Controller_0:avs_s0_read
	signal mm_interconnect_0_ng_controller_0_s0_byteenable                                 : std_logic_vector(3 downto 0);  -- mm_interconnect_0:NG_Controller_0_s0_byteenable -> NG_Controller_0:avs_s0_byteenable
	signal mm_interconnect_0_ng_controller_0_s0_write                                      : std_logic;                     -- mm_interconnect_0:NG_Controller_0_s0_write -> NG_Controller_0:avs_s0_write
	signal mm_interconnect_0_ng_controller_0_s0_writedata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:NG_Controller_0_s0_writedata -> NG_Controller_0:avs_s0_writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect                                : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata                                  : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address                                   : std_logic_vector(9 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable                                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write                                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal irq_mapper_receiver0_irq                                                        : std_logic;                     -- OY_MM_Controller_0:ins_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                        : std_logic;                     -- TEST_OY_Controller_0:ins_irq -> irq_mapper:receiver1_irq
	signal nios2_gen2_0_irq_irq                                                            : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                                                  : std_logic;                     -- rst_controller:reset_out -> [NG_Controller_0:rsi_reset, TEST_OY_Controller_0:rsi_reset, irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                              : std_logic;                     -- rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                                              : std_logic;                     -- rst_controller_001:reset_out -> [OY_MM_Controller_0:rsi_reset, mm_interconnect_0:OY_MM_Controller_0_reset_reset_bridge_in_reset_reset]
	signal rst_controller_reset_out_reset_ports_inv                                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [NG_Instr_Controller_0:resetn, nios2_gen2_0:reset_n]

begin

	ng_controller_0 : component Number_generator_controller
		port map (
			avs_s0_chipselect => mm_interconnect_0_ng_controller_0_s0_chipselect, --    s0.chipselect
			avs_s0_byteenable => mm_interconnect_0_ng_controller_0_s0_byteenable, --      .byteenable
			avs_s0_read       => mm_interconnect_0_ng_controller_0_s0_read,       --      .read
			avs_s0_readdata   => mm_interconnect_0_ng_controller_0_s0_readdata,   --      .readdata
			avs_s0_write      => mm_interconnect_0_ng_controller_0_s0_write,      --      .write
			avs_s0_writedata  => mm_interconnect_0_ng_controller_0_s0_writedata,  --      .writedata
			csi_clk           => clk_clk,                                         -- clock.clk
			rsi_reset         => rst_controller_reset_out_reset                   -- reset.reset
		);

	ng_instr_controller_0 : component CI_NG
		port map (
			clk    => clk_clk,                                                                        --                         clock.clk
			result => nios2_gen2_0_custom_instruction_master_comb_slave_translator0_ci_master_result, -- nios_custom_instruction_slave.result
			resetn => rst_controller_reset_out_reset_ports_inv                                        --                         reset.reset_n
		);

	oy_instr_controller_0 : component OY_Instruction_Controller
		generic map (
			n => 16
		)
		port map (
			ncs_clk    => nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_clk,    -- nios_custom_instruction_slave.clk
			ncs_reset  => nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_reset,  --                              .reset
			ncs_start  => nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_start,  --                              .start
			ncs_dataa  => nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_dataa,  --                              .dataa
			ncs_datab  => nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_datab,  --                              .datab
			ncs_done   => nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_done,   --                              .done
			ncs_result => nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_result  --                              .result
		);

	oy_mm_controller_0 : component OY_MM_Controller
		generic map (
			n => 16
		)
		port map (
			avs_chipselect  => mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_chipselect,  --     avalon_slave_0.chipselect
			avs_address     => mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_address,     --                   .address
			avs_read        => mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_read,        --                   .read
			avs_readdata    => mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_readdata,    --                   .readdata
			avs_write       => mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_write,       --                   .write
			avs_writedata   => mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_writedata,   --                   .writedata
			avs_byteenable  => mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_byteenable,  --                   .byteenable
			avs_waitrequest => mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_waitrequest, --                   .waitrequest
			csi_clk         => clk_clk,                                                         --              clock.clk
			rsi_reset       => rst_controller_001_reset_out_reset,                              --              reset.reset
			ins_irq         => irq_mapper_receiver0_irq                                         -- interrupt_sender_0.irq
		);

	test_oy_controller_0 : component TEST_OY_Controller
		generic map (
			n => 16
		)
		port map (
			avs_chipselect  => mm_interconnect_0_test_oy_controller_0_avalon_slave_0_chipselect,  --     avalon_slave_0.chipselect
			avs_address     => mm_interconnect_0_test_oy_controller_0_avalon_slave_0_address,     --                   .address
			avs_read        => mm_interconnect_0_test_oy_controller_0_avalon_slave_0_read,        --                   .read
			avs_readdata    => mm_interconnect_0_test_oy_controller_0_avalon_slave_0_readdata,    --                   .readdata
			avs_write       => mm_interconnect_0_test_oy_controller_0_avalon_slave_0_write,       --                   .write
			avs_writedata   => mm_interconnect_0_test_oy_controller_0_avalon_slave_0_writedata,   --                   .writedata
			avs_byteenable  => mm_interconnect_0_test_oy_controller_0_avalon_slave_0_byteenable,  --                   .byteenable
			avs_waitrequest => mm_interconnect_0_test_oy_controller_0_avalon_slave_0_waitrequest, --                   .waitrequest
			csi_clk         => clk_clk,                                                           --              clock.clk
			rsi_reset       => rst_controller_reset_out_reset,                                    --              reset.reset
			ins_irq         => irq_mapper_receiver1_irq                                           -- interrupt_sender_0.irq
		);

	nios2_gen2_0 : component TEST_OY_CPU_nios2_gen2_0
		port map (
			clk                                 => clk_clk,                                                    --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                   --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                         --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			E_ci_multi_done                     => nios2_gen2_0_custom_instruction_master_done,                -- custom_instruction_master.done
			E_ci_multi_clk_en                   => nios2_gen2_0_custom_instruction_master_clk_en,              --                          .clk_en
			E_ci_multi_start                    => nios2_gen2_0_custom_instruction_master_start,               --                          .start
			E_ci_result                         => nios2_gen2_0_custom_instruction_master_result,              --                          .result
			D_ci_a                              => nios2_gen2_0_custom_instruction_master_a,                   --                          .a
			D_ci_b                              => nios2_gen2_0_custom_instruction_master_b,                   --                          .b
			D_ci_c                              => nios2_gen2_0_custom_instruction_master_c,                   --                          .c
			D_ci_n                              => nios2_gen2_0_custom_instruction_master_n,                   --                          .n
			D_ci_readra                         => nios2_gen2_0_custom_instruction_master_readra,              --                          .readra
			D_ci_readrb                         => nios2_gen2_0_custom_instruction_master_readrb,              --                          .readrb
			D_ci_writerc                        => nios2_gen2_0_custom_instruction_master_writerc,             --                          .writerc
			E_ci_dataa                          => nios2_gen2_0_custom_instruction_master_dataa,               --                          .dataa
			E_ci_datab                          => nios2_gen2_0_custom_instruction_master_datab,               --                          .datab
			E_ci_multi_clock                    => nios2_gen2_0_custom_instruction_master_clk,                 --                          .clk
			E_ci_multi_reset                    => nios2_gen2_0_custom_instruction_master_reset,               --                          .reset
			E_ci_multi_reset_req                => nios2_gen2_0_custom_instruction_master_reset_req,           --                          .reset_req
			W_ci_estatus                        => nios2_gen2_0_custom_instruction_master_estatus,             --                          .estatus
			W_ci_ipending                       => nios2_gen2_0_custom_instruction_master_ipending             --                          .ipending
		);

	onchip_memory2_0 : component TEST_OY_CPU_onchip_memory2_0
		port map (
			clk        => clk_clk,                                          --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,               --       .reset_req
			freeze     => '0'                                               -- (terminated)
		);

	nios2_gen2_0_custom_instruction_master_translator : component altera_customins_master_translator
		generic map (
			SHARED_COMB_AND_MULTI => 1
		)
		port map (
			ci_slave_dataa            => nios2_gen2_0_custom_instruction_master_dataa,                                --        ci_slave.dataa
			ci_slave_datab            => nios2_gen2_0_custom_instruction_master_datab,                                --                .datab
			ci_slave_result           => nios2_gen2_0_custom_instruction_master_result,                               --                .result
			ci_slave_n                => nios2_gen2_0_custom_instruction_master_n,                                    --                .n
			ci_slave_readra           => nios2_gen2_0_custom_instruction_master_readra,                               --                .readra
			ci_slave_readrb           => nios2_gen2_0_custom_instruction_master_readrb,                               --                .readrb
			ci_slave_writerc          => nios2_gen2_0_custom_instruction_master_writerc,                              --                .writerc
			ci_slave_a                => nios2_gen2_0_custom_instruction_master_a,                                    --                .a
			ci_slave_b                => nios2_gen2_0_custom_instruction_master_b,                                    --                .b
			ci_slave_c                => nios2_gen2_0_custom_instruction_master_c,                                    --                .c
			ci_slave_ipending         => nios2_gen2_0_custom_instruction_master_ipending,                             --                .ipending
			ci_slave_estatus          => nios2_gen2_0_custom_instruction_master_estatus,                              --                .estatus
			ci_slave_multi_clk        => nios2_gen2_0_custom_instruction_master_clk,                                  --                .clk
			ci_slave_multi_reset      => nios2_gen2_0_custom_instruction_master_reset,                                --                .reset
			ci_slave_multi_clken      => nios2_gen2_0_custom_instruction_master_clk_en,                               --                .clk_en
			ci_slave_multi_reset_req  => nios2_gen2_0_custom_instruction_master_reset_req,                            --                .reset_req
			ci_slave_multi_start      => nios2_gen2_0_custom_instruction_master_start,                                --                .start
			ci_slave_multi_done       => nios2_gen2_0_custom_instruction_master_done,                                 --                .done
			comb_ci_master_dataa      => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_dataa,      --  comb_ci_master.dataa
			comb_ci_master_datab      => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_datab,      --                .datab
			comb_ci_master_result     => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_result,     --                .result
			comb_ci_master_n          => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_n,          --                .n
			comb_ci_master_readra     => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_readra,     --                .readra
			comb_ci_master_readrb     => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_readrb,     --                .readrb
			comb_ci_master_writerc    => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_writerc,    --                .writerc
			comb_ci_master_a          => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_a,          --                .a
			comb_ci_master_b          => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_b,          --                .b
			comb_ci_master_c          => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_c,          --                .c
			comb_ci_master_ipending   => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_ipending,   --                .ipending
			comb_ci_master_estatus    => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_estatus,    --                .estatus
			multi_ci_master_clk       => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_clk,       -- multi_ci_master.clk
			multi_ci_master_reset     => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_reset,     --                .reset
			multi_ci_master_clken     => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_clk_en,    --                .clk_en
			multi_ci_master_reset_req => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_reset_req, --                .reset_req
			multi_ci_master_start     => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_start,     --                .start
			multi_ci_master_done      => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_done,      --                .done
			multi_ci_master_dataa     => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_dataa,     --                .dataa
			multi_ci_master_datab     => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_datab,     --                .datab
			multi_ci_master_result    => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_result,    --                .result
			multi_ci_master_n         => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_n,         --                .n
			multi_ci_master_readra    => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_readra,    --                .readra
			multi_ci_master_readrb    => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_readrb,    --                .readrb
			multi_ci_master_writerc   => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_writerc,   --                .writerc
			multi_ci_master_a         => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_a,         --                .a
			multi_ci_master_b         => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_b,         --                .b
			multi_ci_master_c         => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_c,         --                .c
			ci_slave_multi_dataa      => "00000000000000000000000000000000",                                          --     (terminated)
			ci_slave_multi_datab      => "00000000000000000000000000000000",                                          --     (terminated)
			ci_slave_multi_result     => open,                                                                        --     (terminated)
			ci_slave_multi_n          => "00000000",                                                                  --     (terminated)
			ci_slave_multi_readra     => '0',                                                                         --     (terminated)
			ci_slave_multi_readrb     => '0',                                                                         --     (terminated)
			ci_slave_multi_writerc    => '0',                                                                         --     (terminated)
			ci_slave_multi_a          => "00000",                                                                     --     (terminated)
			ci_slave_multi_b          => "00000",                                                                     --     (terminated)
			ci_slave_multi_c          => "00000"                                                                      --     (terminated)
		);

	nios2_gen2_0_custom_instruction_master_comb_xconnect : component TEST_OY_CPU_nios2_gen2_0_custom_instruction_master_comb_xconnect
		port map (
			ci_slave_dataa      => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_dataa,    --   ci_slave.dataa
			ci_slave_datab      => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_datab,    --           .datab
			ci_slave_result     => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_result,   --           .result
			ci_slave_n          => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_n,        --           .n
			ci_slave_readra     => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_readra,   --           .readra
			ci_slave_readrb     => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_readrb,   --           .readrb
			ci_slave_writerc    => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_writerc,  --           .writerc
			ci_slave_a          => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_a,        --           .a
			ci_slave_b          => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_b,        --           .b
			ci_slave_c          => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_c,        --           .c
			ci_slave_ipending   => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_ipending, --           .ipending
			ci_slave_estatus    => nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_estatus,  --           .estatus
			ci_master0_dataa    => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_dataa,     -- ci_master0.dataa
			ci_master0_datab    => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_datab,     --           .datab
			ci_master0_result   => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_result,    --           .result
			ci_master0_n        => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_n,         --           .n
			ci_master0_readra   => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_readra,    --           .readra
			ci_master0_readrb   => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_readrb,    --           .readrb
			ci_master0_writerc  => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_writerc,   --           .writerc
			ci_master0_a        => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_a,         --           .a
			ci_master0_b        => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_b,         --           .b
			ci_master0_c        => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_c,         --           .c
			ci_master0_ipending => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_ipending,  --           .ipending
			ci_master0_estatus  => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_estatus    --           .estatus
		);

	nios2_gen2_0_custom_instruction_master_comb_slave_translator0 : component test_oy_cpu_nios2_gen2_0_custom_instruction_master_comb_slave_translator0
		generic map (
			N_WIDTH          => 8,
			USE_DONE         => 0,
			NUM_FIXED_CYCLES => 0
		)
		port map (
			ci_slave_dataa      => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_dataa,          --  ci_slave.dataa
			ci_slave_datab      => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_datab,          --          .datab
			ci_slave_result     => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_result,         --          .result
			ci_slave_n          => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_n,              --          .n
			ci_slave_readra     => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_readra,         --          .readra
			ci_slave_readrb     => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_readrb,         --          .readrb
			ci_slave_writerc    => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_writerc,        --          .writerc
			ci_slave_a          => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_a,              --          .a
			ci_slave_b          => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_b,              --          .b
			ci_slave_c          => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_c,              --          .c
			ci_slave_ipending   => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_ipending,       --          .ipending
			ci_slave_estatus    => nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_estatus,        --          .estatus
			ci_master_result    => nios2_gen2_0_custom_instruction_master_comb_slave_translator0_ci_master_result, -- ci_master.result
			ci_master_dataa     => open,                                                                           -- (terminated)
			ci_master_datab     => open,                                                                           -- (terminated)
			ci_master_n         => open,                                                                           -- (terminated)
			ci_master_readra    => open,                                                                           -- (terminated)
			ci_master_readrb    => open,                                                                           -- (terminated)
			ci_master_writerc   => open,                                                                           -- (terminated)
			ci_master_a         => open,                                                                           -- (terminated)
			ci_master_b         => open,                                                                           -- (terminated)
			ci_master_c         => open,                                                                           -- (terminated)
			ci_master_ipending  => open,                                                                           -- (terminated)
			ci_master_estatus   => open,                                                                           -- (terminated)
			ci_master_clk       => open,                                                                           -- (terminated)
			ci_master_clken     => open,                                                                           -- (terminated)
			ci_master_reset_req => open,                                                                           -- (terminated)
			ci_master_reset     => open,                                                                           -- (terminated)
			ci_master_start     => open,                                                                           -- (terminated)
			ci_master_done      => '0',                                                                            -- (terminated)
			ci_slave_clk        => '0',                                                                            -- (terminated)
			ci_slave_clken      => '0',                                                                            -- (terminated)
			ci_slave_reset_req  => '0',                                                                            -- (terminated)
			ci_slave_reset      => '0',                                                                            -- (terminated)
			ci_slave_start      => '0',                                                                            -- (terminated)
			ci_slave_done       => open                                                                            -- (terminated)
		);

	nios2_gen2_0_custom_instruction_master_multi_xconnect : component TEST_OY_CPU_nios2_gen2_0_custom_instruction_master_multi_xconnect
		port map (
			ci_slave_dataa       => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_dataa,     --   ci_slave.dataa
			ci_slave_datab       => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_datab,     --           .datab
			ci_slave_result      => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_result,    --           .result
			ci_slave_n           => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_n,         --           .n
			ci_slave_readra      => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_readra,    --           .readra
			ci_slave_readrb      => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_readrb,    --           .readrb
			ci_slave_writerc     => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_writerc,   --           .writerc
			ci_slave_a           => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_a,         --           .a
			ci_slave_b           => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_b,         --           .b
			ci_slave_c           => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_c,         --           .c
			ci_slave_ipending    => open,                                                                        --           .ipending
			ci_slave_estatus     => open,                                                                        --           .estatus
			ci_slave_clk         => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_clk,       --           .clk
			ci_slave_reset       => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_reset,     --           .reset
			ci_slave_clken       => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_clk_en,    --           .clk_en
			ci_slave_reset_req   => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_reset_req, --           .reset_req
			ci_slave_start       => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_start,     --           .start
			ci_slave_done        => nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_done,      --           .done
			ci_master0_dataa     => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_dataa,      -- ci_master0.dataa
			ci_master0_datab     => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_datab,      --           .datab
			ci_master0_result    => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_result,     --           .result
			ci_master0_n         => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_n,          --           .n
			ci_master0_readra    => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_readra,     --           .readra
			ci_master0_readrb    => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_readrb,     --           .readrb
			ci_master0_writerc   => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_writerc,    --           .writerc
			ci_master0_a         => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_a,          --           .a
			ci_master0_b         => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_b,          --           .b
			ci_master0_c         => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_c,          --           .c
			ci_master0_ipending  => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_ipending,   --           .ipending
			ci_master0_estatus   => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_estatus,    --           .estatus
			ci_master0_clk       => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_clk,        --           .clk
			ci_master0_reset     => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_reset,      --           .reset
			ci_master0_clken     => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_clk_en,     --           .clk_en
			ci_master0_reset_req => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_reset_req,  --           .reset_req
			ci_master0_start     => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_start,      --           .start
			ci_master0_done      => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_done        --           .done
		);

	nios2_gen2_0_custom_instruction_master_multi_slave_translator0 : component test_oy_cpu_nios2_gen2_0_custom_instruction_master_multi_slave_translator0
		generic map (
			N_WIDTH          => 8,
			USE_DONE         => 1,
			NUM_FIXED_CYCLES => 0
		)
		port map (
			ci_slave_dataa      => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_dataa,          --  ci_slave.dataa
			ci_slave_datab      => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_datab,          --          .datab
			ci_slave_result     => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_result,         --          .result
			ci_slave_n          => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_n,              --          .n
			ci_slave_readra     => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_readra,         --          .readra
			ci_slave_readrb     => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_readrb,         --          .readrb
			ci_slave_writerc    => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_writerc,        --          .writerc
			ci_slave_a          => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_a,              --          .a
			ci_slave_b          => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_b,              --          .b
			ci_slave_c          => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_c,              --          .c
			ci_slave_ipending   => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_ipending,       --          .ipending
			ci_slave_estatus    => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_estatus,        --          .estatus
			ci_slave_clk        => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_clk,            --          .clk
			ci_slave_clken      => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_clk_en,         --          .clk_en
			ci_slave_reset_req  => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_reset_req,      --          .reset_req
			ci_slave_reset      => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_reset,          --          .reset
			ci_slave_start      => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_start,          --          .start
			ci_slave_done       => nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_done,           --          .done
			ci_master_dataa     => nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_dataa,  -- ci_master.dataa
			ci_master_datab     => nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_datab,  --          .datab
			ci_master_result    => nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_result, --          .result
			ci_master_clk       => nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_clk,    --          .clk
			ci_master_clken     => open,                                                                            --          .clk_en
			ci_master_reset     => nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_reset,  --          .reset
			ci_master_start     => nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_start,  --          .start
			ci_master_done      => nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_done,   --          .done
			ci_master_n         => open,                                                                            -- (terminated)
			ci_master_readra    => open,                                                                            -- (terminated)
			ci_master_readrb    => open,                                                                            -- (terminated)
			ci_master_writerc   => open,                                                                            -- (terminated)
			ci_master_a         => open,                                                                            -- (terminated)
			ci_master_b         => open,                                                                            -- (terminated)
			ci_master_c         => open,                                                                            -- (terminated)
			ci_master_ipending  => open,                                                                            -- (terminated)
			ci_master_estatus   => open,                                                                            -- (terminated)
			ci_master_reset_req => open                                                                             -- (terminated)
		);

	mm_interconnect_0 : component TEST_OY_CPU_mm_interconnect_0
		port map (
			clk_0_clk_clk                                        => clk_clk,                                                           --                                      clk_0_clk.clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset       => rst_controller_reset_out_reset,                                    --       nios2_gen2_0_reset_reset_bridge_in_reset.reset
			OY_MM_Controller_0_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                                -- OY_MM_Controller_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address                     => nios2_gen2_0_data_master_address,                                  --                       nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest                 => nios2_gen2_0_data_master_waitrequest,                              --                                               .waitrequest
			nios2_gen2_0_data_master_byteenable                  => nios2_gen2_0_data_master_byteenable,                               --                                               .byteenable
			nios2_gen2_0_data_master_read                        => nios2_gen2_0_data_master_read,                                     --                                               .read
			nios2_gen2_0_data_master_readdata                    => nios2_gen2_0_data_master_readdata,                                 --                                               .readdata
			nios2_gen2_0_data_master_write                       => nios2_gen2_0_data_master_write,                                    --                                               .write
			nios2_gen2_0_data_master_writedata                   => nios2_gen2_0_data_master_writedata,                                --                                               .writedata
			nios2_gen2_0_data_master_debugaccess                 => nios2_gen2_0_data_master_debugaccess,                              --                                               .debugaccess
			nios2_gen2_0_instruction_master_address              => nios2_gen2_0_instruction_master_address,                           --                nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest          => nios2_gen2_0_instruction_master_waitrequest,                       --                                               .waitrequest
			nios2_gen2_0_instruction_master_read                 => nios2_gen2_0_instruction_master_read,                              --                                               .read
			nios2_gen2_0_instruction_master_readdata             => nios2_gen2_0_instruction_master_readdata,                          --                                               .readdata
			NG_Controller_0_s0_write                             => mm_interconnect_0_ng_controller_0_s0_write,                        --                             NG_Controller_0_s0.write
			NG_Controller_0_s0_read                              => mm_interconnect_0_ng_controller_0_s0_read,                         --                                               .read
			NG_Controller_0_s0_readdata                          => mm_interconnect_0_ng_controller_0_s0_readdata,                     --                                               .readdata
			NG_Controller_0_s0_writedata                         => mm_interconnect_0_ng_controller_0_s0_writedata,                    --                                               .writedata
			NG_Controller_0_s0_byteenable                        => mm_interconnect_0_ng_controller_0_s0_byteenable,                   --                                               .byteenable
			NG_Controller_0_s0_chipselect                        => mm_interconnect_0_ng_controller_0_s0_chipselect,                   --                                               .chipselect
			nios2_gen2_0_debug_mem_slave_address                 => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,            --                   nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write                   => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,              --                                               .write
			nios2_gen2_0_debug_mem_slave_read                    => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,               --                                               .read
			nios2_gen2_0_debug_mem_slave_readdata                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,           --                                               .readdata
			nios2_gen2_0_debug_mem_slave_writedata               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,          --                                               .writedata
			nios2_gen2_0_debug_mem_slave_byteenable              => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,         --                                               .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,        --                                               .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,        --                                               .debugaccess
			onchip_memory2_0_s1_address                          => mm_interconnect_0_onchip_memory2_0_s1_address,                     --                            onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                            => mm_interconnect_0_onchip_memory2_0_s1_write,                       --                                               .write
			onchip_memory2_0_s1_readdata                         => mm_interconnect_0_onchip_memory2_0_s1_readdata,                    --                                               .readdata
			onchip_memory2_0_s1_writedata                        => mm_interconnect_0_onchip_memory2_0_s1_writedata,                   --                                               .writedata
			onchip_memory2_0_s1_byteenable                       => mm_interconnect_0_onchip_memory2_0_s1_byteenable,                  --                                               .byteenable
			onchip_memory2_0_s1_chipselect                       => mm_interconnect_0_onchip_memory2_0_s1_chipselect,                  --                                               .chipselect
			onchip_memory2_0_s1_clken                            => mm_interconnect_0_onchip_memory2_0_s1_clken,                       --                                               .clken
			OY_MM_Controller_0_avalon_slave_0_address            => mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_address,       --              OY_MM_Controller_0_avalon_slave_0.address
			OY_MM_Controller_0_avalon_slave_0_write              => mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_write,         --                                               .write
			OY_MM_Controller_0_avalon_slave_0_read               => mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_read,          --                                               .read
			OY_MM_Controller_0_avalon_slave_0_readdata           => mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_readdata,      --                                               .readdata
			OY_MM_Controller_0_avalon_slave_0_writedata          => mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_writedata,     --                                               .writedata
			OY_MM_Controller_0_avalon_slave_0_byteenable         => mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_byteenable,    --                                               .byteenable
			OY_MM_Controller_0_avalon_slave_0_waitrequest        => mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_waitrequest,   --                                               .waitrequest
			OY_MM_Controller_0_avalon_slave_0_chipselect         => mm_interconnect_0_oy_mm_controller_0_avalon_slave_0_chipselect,    --                                               .chipselect
			TEST_OY_Controller_0_avalon_slave_0_address          => mm_interconnect_0_test_oy_controller_0_avalon_slave_0_address,     --            TEST_OY_Controller_0_avalon_slave_0.address
			TEST_OY_Controller_0_avalon_slave_0_write            => mm_interconnect_0_test_oy_controller_0_avalon_slave_0_write,       --                                               .write
			TEST_OY_Controller_0_avalon_slave_0_read             => mm_interconnect_0_test_oy_controller_0_avalon_slave_0_read,        --                                               .read
			TEST_OY_Controller_0_avalon_slave_0_readdata         => mm_interconnect_0_test_oy_controller_0_avalon_slave_0_readdata,    --                                               .readdata
			TEST_OY_Controller_0_avalon_slave_0_writedata        => mm_interconnect_0_test_oy_controller_0_avalon_slave_0_writedata,   --                                               .writedata
			TEST_OY_Controller_0_avalon_slave_0_byteenable       => mm_interconnect_0_test_oy_controller_0_avalon_slave_0_byteenable,  --                                               .byteenable
			TEST_OY_Controller_0_avalon_slave_0_waitrequest      => mm_interconnect_0_test_oy_controller_0_avalon_slave_0_waitrequest, --                                               .waitrequest
			TEST_OY_Controller_0_avalon_slave_0_chipselect       => mm_interconnect_0_test_oy_controller_0_avalon_slave_0_chipselect   --                                               .chipselect
		);

	irq_mapper : component TEST_OY_CPU_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => nios2_gen2_0_irq_irq            --    sender.irq
		);

	rst_controller : component test_oy_cpu_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_gen2_0_debug_reset_request_reset, -- reset_in0.reset
			reset_in1      => nios2_gen2_0_debug_reset_request_reset, -- reset_in1.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_reset_out_reset,         -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,     --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_001 : component test_oy_cpu_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_gen2_0_debug_reset_request_reset, -- reset_in0.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => open,                                   -- (terminated)
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of TEST_OY_CPU
